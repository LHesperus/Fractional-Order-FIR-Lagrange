library verilog;
use verilog.vl_types.all;
entity int_delay_tb is
end int_delay_tb;
